parameter TX_SIZE = 1024;